//=============================================================================
// Project  : HoneyB V2
// File Name: xlr_gpp_pkg.sv
//=============================================================================
// Description: Package for agent xlr_gpp
//=============================================================================

package xlr_gpp_pkg;

// Empty package

endpackage : xlr_gpp_pkg
