//=============================================================================
// Project  : HoneyB V2
// File Name: top_pkg.sv
//=============================================================================
// Description: Package for top
//=============================================================================

package top_pkg;

//  `include "uvm_macros.svh"

//  import uvm_pkg::*;

//  import xlr_mem_pkg::*;
//  import xlr_gpp_pkg::*;

//  `include "top_config.sv"
//  `include "top_seq_lib.sv"
//  `include "port_converter.sv"
//  `include "reference.sv"
//  `include "top_env.sv"
//  `include "xlr_scoreboard.sv"

endpackage : top_pkg

