//=========================================================================================
// Project  : HoneyB V1
// File Name: xlr_mem_monitor.sv
//=========================================================================================
// Description: Monitor for xlr_mem
// Important: The monitor takes care both of the inputs and the outputs
//            therefore it has 2 analysis ports, 1 for the inputs and 1 for outputs
//            since we have a single tx class for both input & output
//            this means that the transaction being broadcasted includes all tx's
//            thus, through the input analysis ports the output signals will be
//            propagated with 'x' values and vice versa for the output analysis port.
//=========================================================================================

`ifndef XLR_MEM_MONITOR_SV
`define XLR_MEM_MONITOR_SV

`include "uvm_macros.svh"
import uvm_pkg::*;
import honeyb_pkg::*;

class xlr_mem_monitor extends uvm_monitor;

  `uvm_component_utils(xlr_mem_monitor)

  virtual xlr_mem_if vif;

  uvm_analysis_port #(xlr_mem_tx) analysis_port_in; // input signals
  uvm_analysis_port #(xlr_mem_tx) analysis_port_out; // output signals

  xlr_mem_tx m_trans_in;
  xlr_mem_tx m_trans_out;

  extern function new(string name, uvm_component parent);

  // Methods build_phase, run_phase, and do_mon generated by setting monitor_inc in file xlr_mem.tpl
  extern function void build_phase(uvm_phase phase);
  extern task run_phase(uvm_phase phase);
  extern task do_mon();
endclass : xlr_mem_monitor 


function xlr_mem_monitor::new(string name, uvm_component parent);
  super.new(name, parent);
  analysis_port_in = new("analysis_port_in", this);
  analysis_port_out = new("analysis_port_out", this);
endfunction : new


function void xlr_mem_monitor::build_phase(uvm_phase phase);
endfunction : build_phase


task xlr_mem_monitor::run_phase(uvm_phase phase);
  `uvm_info("", "run_phase", UVM_NONE)
  m_trans_in = xlr_mem_tx::type_id::create("m_trans_in");
  m_trans_out = xlr_mem_tx::type_id::create("m_trans_out");
  do_mon();
endtask : run_phase

task xlr_mem_monitor::do_mon();

  bit rd_sent = 1'b0; // Flag for read request
  bit wr_sent = 1'b0; // Flag for write request
  bit rst_asserted = 1'b0; // Flag for rst_n
  bit first_rd = 1'b1; // a stupid implementation to get rid of annoying msg I don't have the patience to deal with
  bit first_wr = 1'b1; // same

  fork // in / out monitors work in parallel

    //*********************************************************************//
    //                           DUT INPUT MONITOR                         //
    //---------------------------------------------------------------------//
    //     Monitor only when in reg's asserted (indicating valid input)    //
    //     Inputs are testbench related (by driver) and set to be sent on  //
    //     negedge Making sure that no timing violations will occur        //
    //                                                                     //
    //*********************************************************************//

    // Input rst_n handling.
    forever begin
      if (!vif.rst_n) begin
        rst_asserted = 1'b1;
        #1; // add small delay
        m_trans_in.mem_rdata = '0;
        `honeyb("MEM MON", "rst_n detected, INPUT transactions are reset")
        analysis_port_in.write(m_trans_in);
      end
      @(vif.rst_n); // Wait until rst_n changes.
      rst_asserted = 1'b0;
    end

    forever @(negedge vif.clk) begin
      #1; // small delay so it can capture the driver's NBA assignments.
      // Always Capture the input values
      m_trans_in.mem_rdata = vif.mem_rdata;

      // If statements to decide when to broadcast and where
      if (vif.mem_rd == 1'b1) begin // optional - add the addr[0] == '0; if we want
        m_trans_in.mem_rd = vif.mem_rd; // pass it through the transaction for REF Model - Important
        m_trans_in.mem_addr = vif.mem_addr; // pass it for REF too.
        // Log the captured data
        `uvm_info("MEM MON", $sformatf("\nRead Requested! Addr SRC : mem_addr[0] = %0d", vif.mem_addr[0]), UVM_MEDIUM);
        `uvm_info("MEM MON", $sformatf("\nmem_rdata[0][0] = %0d\nmem_rdata[0][1] = %0d\nmem_rdata[0][2]] = %0d\nmem_rdata[0][3] = %0d\nmem_rdata[0][4] = %0d\nmem_rdata[0][5] = %0d\nmem_rdata[0][6] = %0d\nmem_rdata[0][7] = %0d", m_trans_in.mem_rdata[0][0], m_trans_in.mem_rdata[0][1], m_trans_in.mem_rdata[0][2], m_trans_in.mem_rdata[0][3], m_trans_in.mem_rdata[0][4], m_trans_in.mem_rdata[0][5], m_trans_in.mem_rdata[0][6], m_trans_in.mem_rdata[0][7]), UVM_MEDIUM);
        rd_sent = 1'b1; // Set rd_sent
        wr_sent = 1'b0; // Reset wr_sent
        first_rd = 1'b0;
        analysis_port_in.write(m_trans_in); // broadcast to REF
      end
    end

    //*********************************************************************//
    //                           DUT OUTPUT MONITOR                        //
    //---------------------------------------------------------------------//
    //     Monitor only when out reg's asserted (indicating valid output)  //
    //     Outputs are DUT related and set to be sent on posedge.          //
    //     This will allow well synchronized timing of the triggerd        //
    //     signals from the DUT.                                           //
    //                                                                     //
    //*********************************************************************//

    // Output rst_n handling.
    forever begin
      if (!vif.rst_n) begin
        #1;
        m_trans_out.mem_addr = vif.mem_addr;
        m_trans_out.mem_wdata = vif.mem_wdata;
        m_trans_out.mem_be = vif.mem_be;
        m_trans_out.mem_rd = vif.mem_rd;
        m_trans_out.mem_wr = vif.mem_wr;
        `uvm_info("MEM MON", "\nrst_n detected, expecting DUT to drive zero OUTPUTS", UVM_MEDIUM);
        analysis_port_out.write(m_trans_out);
      end
      @(vif.rst_n); // Wait until rst_n changes.
    end

    forever @(posedge vif.clk) begin
      // Always capture the output values
      m_trans_out.mem_addr = vif.mem_addr;
      m_trans_out.mem_wdata = vif.mem_wdata;
      m_trans_out.mem_be = vif.mem_be;
      m_trans_out.mem_rd = vif.mem_rd;
      m_trans_out.mem_wr = vif.mem_wr;

      // If statements to decide if, when & where to broadcast
      if (vif.mem_wr == 1'b1) begin
        // Log the captured data
        `uvm_info("MEM MON", $sformatf("\nWrite Requested! Addr SRC : mem_addr[0] = %0d", m_trans_out.mem_addr[0]), UVM_MEDIUM);
        wr_sent = 1'b1; // Set wr_sent
        rd_sent = 1'b0; // Reset rd_sent
        first_wr = 1'b0;
        analysis_port_out.write(m_trans_out); // Broadcast to scoreboard
      end
    end
  join
endtask : do_mon

`endif // XLR_MEM_MONITOR_SV

