//=========================================================================================
// Project  : HoneyB V2
// File Name: xlr_mem_monitor.sv
//=========================================================================================
// Description: Monitor for xlr_mem
// Important: The monitor takes care both of the inputs and the outputs
//            therefore it has 2 analysis ports, 1 for the inputs and 1 for outputs
//            since we have a single tx class for both input & output
//            this means that the transaction being broadcasted includes all tx's
//            thus, through the input analysis ports the output signals will be
//            propagated with 'x' values and vice versa for the output analysis port.
//=========================================================================================

`ifndef XLR_MEM_MONITOR_SV
`define XLR_MEM_MONITOR_SV

`include "uvm_macros.svh"
import uvm_pkg::*;
import honeyb_pkg::*;
import xlr_mem_pkg::*;

class xlr_mem_monitor extends uvm_monitor;

    `uvm_component_utils(xlr_mem_monitor)

    /* Monitor accesses parameterized interface through a reference to the abstract base class
      NOTE - Even though importing the pkg, I use it this way to emphasize the change, may simplify later*/

    virtual xlr_mem_if vif; // OLD
    xlr_mem_pkg::xlr_mem_if_base m_xlr_mem_if; // NEW

    uvm_analysis_port #(xlr_mem_tx) analysis_port_in; // input signals
    uvm_analysis_port #(xlr_mem_tx) analysis_port_out; // output signals

    xlr_mem_tx m_trans_in;
    xlr_mem_tx m_trans_out;

    extern function new(string name, uvm_component parent);

    // Methods build_phase, run_phase, and do_mon generated by setting monitor_inc in file xlr_mem.tpl
    extern function void build_phase(uvm_phase phase);
    extern task run_phase(uvm_phase phase);
    extern task do_mon();
endclass : xlr_mem_monitor 


function xlr_mem_monitor::new(string name, uvm_component parent);
    super.new(name, parent);
    analysis_port_in = new("analysis_port_in", this);
    analysis_port_out = new("analysis_port_out", this);
endfunction : new


function void xlr_mem_monitor::build_phase(uvm_phase phase);
endfunction : build_phase


task xlr_mem_monitor::run_phase(uvm_phase phase);
    `honeyb("MEM MON", "run_phase initialized...")
    m_trans_in = xlr_mem_tx::type_id::create("m_trans_in");
    m_trans_out = xlr_mem_tx::type_id::create("m_trans_out");
    do_mon();
endtask : run_phase

task xlr_mem_monitor::do_mon();

    bit rd_sent = 1'b0; // Flag for read request
    bit wr_sent = 1'b0; // Flag for write request
    bit rst_asserted = 1'b0; // Flag for rst_n
    bit first_rd = 1'b1; // a stupid implementation to get rid of annoying msg I don't have the patience to deal with
    bit first_wr = 1'b1; // same

    fork // in / out monitors work in parallel

        /*                           DUT INPUT MONITOR                         
            //---------------------------------------------------------------------//
            //     Monitor only when in reg's asserted (indicating valid input)    //
            //     Inputs are testbench related (by driver) and set to be sent on  //
            //     negedge Making sure that no timing violations will occur        //
            //                                                                     //
            //---------------------------------------------------------------------*/

        // Input rst_n handling.
        forever begin
            // if (!vif.rst_n) begin // OLD
            if (!m_xlr_mem_if.get_rst()) begin // NEW
                rst_asserted = 1'b1;
                #1; // add small delay
                m_trans_in.mem_rdata[MEM0] = '0;
                `honeyb("MEM MON", "rst_n detected, INPUT transactions are reset")
                analysis_port_in.write(m_trans_in);
            end
            // @(vif.rst_n); // Wait until rst_n changes || OLD
            m_xlr_mem_if.wait4rst_n(); // Wait until rst_n changes || NEW
            rst_asserted = 1'b0;
        end

        // forever @(negedge vif.clk) begin // OLD
        forever begin // NEW
            m_xlr_mem_if.negedge_clk();
            #1; // small delay so it can capture the driver's NBA assignments.
            // Always Capture the input values
            // m_trans_in.mem_rdata = vif.mem_rdata; // OLD
            m_trans_in.mem_rdata = m_xlr_mem_if.get_mem_rdata(MEM0);
            // If statements to decide when to broadcast and where
            // if (vif.mem_rd == 1'b1) begin // optional - add the addr[0] == '0; if we want || OLD
            if (m_xlr_mem_if.get_mem_rd(MEM0) == 1'b1) begin // optional - add the addr[0] == '0; if we want || NEW
                // m_trans_in.mem_rd = vif.mem_rd; // pass it through the transaction for REF Model - Important || OLD
                m_trans_in.mem_rd[MEM0] = m_xlr_mem_if.get_mem_rd(MEM0); // pass it through the transaction for REF Model - Important || NEW
                // m_trans_in.mem_addr = vif.mem_addr; // pass it for REF too. || OLD
                m_trans_in.mem_addr[MEM0] = m_xlr_mem_if.get_mem_addr(MEM0); // pass it for REF too. || NEW
                // m_trans_in.mem_be = vif.mem_be; // OLD
                m_trans_in.mem_be[MEM0] = m_xlr_mem_if.get_mem_be(MEM0); // NEW
                // Log the captured data
                `honeyb("MEM MON", "Read Requested...")
                m_trans_in.set_mem(MEM0);
                m_trans_in.set_mode("rd");
                m_trans_in.print();
                rd_sent = 1'b1; // Set rd_sent
                wr_sent = 1'b0; // Reset wr_sent
                first_rd = 1'b0;
                analysis_port_in.write(m_trans_in); // broadcast to REF
            end
        end

        /*                           DUT OUTPUT MONITOR                        
            //---------------------------------------------------------------------//
            //     Monitor only when out reg's asserted (indicating valid output)  //
            //     Outputs are DUT related and set to be sent on posedge.          //
            //     This will allow well synchronized timing of the triggerd        //
            //     signals from the DUT.                                           //
            //                                                                     //
            //---------------------------------------------------------------------*/

        // Output rst_n handling.
        forever begin
            // if (!vif.rst_n) begin // OLD
            if (!m_xlr_mem_if.get_rst()) begin // NEW
                #1;
                // m_trans_out.mem_addr = vif.mem_addr; // OLD
                m_trans_out.mem_addr[MEM0] = m_xlr_mem_if.get_mem_addr(MEM0); // NEW

                // m_trans_out.mem_wdata = vif.mem_wdata; // OLD
                m_trans_out.mem_wdata[MEM0] = m_xlr_mem_if.get_mem_wdata(MEM0); // NEW

                // m_trans_out.mem_be = vif.mem_be; // OLD
                m_trans_out.mem_be[MEM0] = m_xlr_mem_if.get_mem_be(MEM0); // NEW

                // m_trans_out.mem_rd = vif.mem_rd; // OLD
                m_trans_out.mem_rd[MEM0] = m_xlr_mem_if.get_mem_rd(MEM0); // NEW

                // m_trans_out.mem_wr = vif.mem_wr; // OLD
                m_trans_out.mem_wr[MEM0] = m_xlr_mem_if.get_mem_wr(MEM0); // NEW
                `honeyb("MEM MON", "rst_n detected, OUTPUT transactions are reset")
                analysis_port_out.write(m_trans_out);
            end
            // @(vif.rst_n); // Wait until rst_n changes || OLD
            m_xlr_mem_if.wait4rst_n(); // Wait until rst_n changes || NEW
        end

        // forever @(posedge vif.clk) begin // OLD
        forever begin // NEW
            m_xlr_mem_if.posedge_clk();
            // Always capture the output values
            // m_trans_out.mem_addr = vif.mem_addr; // OLD
            m_trans_out.mem_addr[MEM0] = m_xlr_mem_if.get_mem_addr(MEM0); // NEW

            // m_trans_out.mem_wdata = vif.mem_wdata; // OLD
            m_trans_out.mem_wdata[MEM0] = m_xlr_mem_if.get_mem_wdata(MEM0); // NEW

            // m_trans_out.mem_be = vif.mem_be; // OLD
            m_trans_out.mem_be[MEM0] = m_xlr_mem_if.get_mem_be(MEM0); // NEW

            // m_trans_out.mem_rd = vif.mem_rd; // OLD
            m_trans_out.mem_rd[MEM0] = m_xlr_mem_if.get_mem_rd(MEM0); // NEW

            // m_trans_out.mem_wr = vif.mem_wr; // OLD
            m_trans_out.mem_wr[MEM0] = m_xlr_mem_if.get_mem_wr(MEM0); // NEW

            // If statements to decide if, when & where to broadcast
            // if (vif.mem_wr == 1'b1) begin // OLD
            if (m_xlr_mem_if.get_mem_wr(MEM0) == 1'b1) begin // NEW
                // Log the captured data
                `honeyb("MEM MON", "Write Requested, Broadcasting...")
                wr_sent = 1'b1; // Set wr_sent
                rd_sent = 1'b0; // Reset rd_sent
                first_wr = 1'b0;
                analysis_port_out.write(m_trans_out); // Broadcast to scoreboard
            end
        end
    join
endtask : do_mon

`endif // XLR_MEM_MONITOR_SV

