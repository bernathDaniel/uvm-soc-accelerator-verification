//=============================================================================
// Project  : HoneyB V1
// File Name: xlr_mem_pkg.sv
//=============================================================================
// Description: Package for agent xlr_mem
//=============================================================================

package xlr_mem_pkg;

// Empty pkg

endpackage : xlr_mem_pkg
