extern function void send_xlr_mem_input(xlr_mem_tx t);
extern function void send_xlr_gpp_input(xlr_gpp_tx t);