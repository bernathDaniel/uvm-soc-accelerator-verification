





    // START CHECK

$monitor("[XLR DUT]: start_honey = %h at %0t", start_honey, $time);  // prints on signal changes
$monitor("[XLR DUT]: xlr_mem_rdata[0] = %h at %0t", xlr_mem_rdata[0], $time);  // prints on signal changes

    // 
